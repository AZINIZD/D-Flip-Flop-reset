//D flip-flop with asynchronous reset (asserted negative)

module dff_reset(D, Clock, Resetn, Q);
    input D, Clock, Resetn;
    output Q;
    reg Q;
 
    always @(negedge Resetn or posedge Clock)
	    if (!Resetn)
            Q <= 0;
        else
            Q <= D;
	
endmodule
